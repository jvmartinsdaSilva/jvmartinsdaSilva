<svg version="1.0" xmlns="http://www.w3.org/2000/svg"
 width="100.000000pt" height="100.000000pt" viewBox="0 0 512.000000 512.000000"
 preserveAspectRatio="xMidYMid meet">

<g transform="translate(0.000000,512.000000) scale(0.100000,-0.100000)"
fill="#ffffff" stroke="none">
<path d="M470 4424 c-221 -47 -408 -236 -455 -459 -22 -105 -22 -2705 0 -2810
47 -225 235 -413 460 -460 105 -22 4065 -22 4170 0 225 47 413 235 460 460 22
105 22 2705 0 2810 -47 225 -235 413 -460 460 -102 21 -4075 21 -4175 -1z
m3989 -402 c-13 -11 -446 -332 -961 -716 l-938 -697 -937 697 c-516 384 -949
705 -962 716 -23 17 30 18 1899 18 1869 0 1922 -1 1899 -18z m-2974 -1112
l1075 -799 1075 799 c591 440 1077 800 1080 800 3 0 4 -562 3 -1248 l-3 -1249
-27 -39 c-15 -21 -44 -50 -65 -64 l-37 -25 -2026 0 -2026 0 -37 25 c-21 14
-50 43 -65 64 l-27 39 -3 1249 c-1 686 0 1248 3 1248 3 0 489 -360 1080 -800z"/>
</g>
</svg>
